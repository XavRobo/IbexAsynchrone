package alu_pkg;

typedef enum logic [4:0] {
ADD,
SUB,
XOR,
OR,
AND,
SRA,
SRL,
SLL,
LT,
LTU,
GE,
GEU,
EQ,
NE,
SLT,
SLTU,
} alu_op;
