//define constqnt used in core

package pkg;

endpackage
