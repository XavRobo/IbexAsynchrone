module tbench_issue;

  //ALU

  logic		     req_alu_o;
  logic [31:0] operand_alu_a;
  logic [31:0] operand_alu_b;
  pkg::alu_op  operateur_alu;

  //pc ALU

  logic [31:0] operand_pc_alu_a;
  logic [31:0] operand_pc_alu_b;
  logic 		   branch_bool;

  //LSU

  logic              data_req;
  logic              data_we;
  logic [31:0]			 lsu_wdata;

  //RF write

  logic [4:0] rf_waddr;
  logic 	    rf_soursel;
  logic 	    req_rf_w;

  issue issue_m (
    .req_i            (req),
    .rst_ni           (rst_ni),
    .rf_rdata_a_i     (rf_rdata_a),
    .rf_rdata_b_i     (rf_rdata_b),
    .pc_rdata_i       (pc_rdata),
    .imm_i_type_i     (imm_i_type),
    .imm_s_type_i     (imm_s_type),
    .imm_b_type_i     (imm_b_type),
    .imm_u_type_i     (imm_u_type),
    .imm_j_type_i     (imm_j_type),
    .imm_o_type_i     (imm_o_type),
    .imm_n_type_i     (imm_n_type),
    .type_operand_a_i (type_operand_a),
    .type_operand_b_i (type_operand_b),
    .type_imm_b_i     (type_imm_b),
    .req_alu_i        (req_alu_o),
    .req_alu_o        (re)
    .operateur_alu_i
  )

endmodule
